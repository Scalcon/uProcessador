library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROM is
	port(	clk     : in std_logic;
			address : in unsigned(6 downto 0);
			instout  : out unsigned(15 downto 0)
		);
end entity;

architecture a_ROM of ROM is
	type mem is array (0 to 127) of unsigned (15 downto 0);
	constant conteudo_rom : mem :=( 
     0 => B"00011111_110_1_1110",
     1 => B"00100000_100_1_1110",
     2 => B"00000010_000_1_1110",
     3 => B"00000010_000_0_1110",
     4 => B"00000000_000_0_1010",
     5 => B"00000000_000_0_0110",
     6 => B"00000001_000_0_1110",
     7 => B"000000000_000_0001",
     8 => B"00000000_000_1_1010",
     9 => B"00000000_000_0_0110",
     10 => B"00000000_110_0_1010",
     11 => B"000000000_000_1100",
     12 => B"00000000_101_1_1010",
     13 => B"00000000_101_0_1010",
     14 => B"000000000_100_0111",
     15 => B"10010_1110101_1101", 
     16 => B"00000000_010_1_1110",
     17 => B"00000010_001_1_1110",
     18 => B"00000010_000_0_1110",
     19 => B"000000000_001_0001",
     20 => B"00000000_001_1_1010",
     21 => B"00000000_010_0_1010",
     22 => B"00000000_001_0_0110",
     23 => B"00000000_110_0_1010",
     24 => B"000000000_001_1100",
     25 => B"00000000_101_1_1010",
     26 => B"00000000_101_0_1010",
     27 => B"000000000_100_0111",
     28 => B"10010_1110110_1101",
     29 => B"00000000_010_1_1110",
     30 => B"00000011_001_1_1110",
     31 => B"00000011_000_0_1110",
     32 => B"000000000_001_0001",
     33 => B"00000000_001_1_1010",
     34 => B"00000000_010_0_1010",
     35 => B"00000000_001_0_0110",
     36 => B"00000000_110_0_1010",
     37 => B"000000000_001_1100",
     38 => B"00000000_101_1_1010",
     39 => B"00000000_101_0_1010",
     40 => B"000000000_100_0111",
     41 => B"10010_1110110_1101",
     42 => B"00000000_010_1_1110",
     43 => B"00000101_001_1_1110",
     44 => B"00000101_000_0_1110",
     45 => B"000000000_001_0001",
     46 => B"00000000_001_1_1010",
     47 => B"00000000_010_0_1010",
     48 => B"00000000_001_0_0110",
     49 => B"00000000_110_0_1010",
     50 => B"000000000_001_1100",
     51 => B"00000000_101_1_1010",
     52 => B"00000000_101_0_1010",
     53 => B"000000000_100_0111",
     54 => B"10010_1110110_1101",
     55 => B"00000000_010_1_1110",
     56 => B"00000111_001_1_1110",
     57 => B"00000111_000_0_1110",
     58 => B"000000000_001_0001",
     59 => B"00000000_001_1_1010",
     60 => B"00000000_010_0_1010",
     61 => B"00000000_001_0_0110",
     62 => B"00000000_110_0_1010",
     63 => B"000000000_001_1100",
     64 => B"00000000_101_1_1010",
     65 => B"00000000_101_0_1010",
     66 => B"000000000_100_0111",
     67 => B"10010_1110110_1101",
     68 => B"00000000_010_1_1110",
     69 => B"00001011_001_1_1110",
     70 => B"00001011_000_0_1110",
     71 => B"000000000_001_0001",
     72 => B"00000000_001_1_1010",
     73 => B"00000000_010_0_1010",
     74 => B"00000000_001_0_0110",
     75 => B"00000000_110_0_1010",
     76 => B"000000000_001_1100",
     77 => B"00000000_101_1_1010",
     78 => B"00000000_101_0_1010",
     79 => B"000000000_100_0111",
     80 => B"10010_1110110_1101",
     81 => B"00000001_000_1_1110",
     82 => B"00000001_000_0_1110",
     83 => B"000000000_000_0001",
     84 => B"00000000_000_1_1010",
     85 => B"00000000_000_1_0110",
     86 => B"00000000_111_1_1010",
     87 => B"00000000_000_0_1010",
     88 => B"000000000_100_0111",
     89 => B"10010_1111001_1101",

		others => (others => '0')
	);
	begin
		
	process(clk) begin
			
		if(rising_edge(clk)) then
			instout <= conteudo_rom(to_integer(address));
		end if;
	end process;
end architecture;	