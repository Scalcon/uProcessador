library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROM is
	port(	clk     : in std_logic;
			address : in unsigned(6 downto 0);
			instout  : out unsigned(15 downto 0)
		);
end entity;

architecture a_ROM of ROM is
	type mem is array (0 to 127) of unsigned (15 downto 0);
	constant conteudo_rom : mem :=( 
     0 => B"00011111_110_1_1110",
     1 => B"00000010_000_1_1110",
     2 => B"00000010_000_0_1110",
     3 => B"00000000_000_0_1010",
     4 => B"00000000_000_0_0110",
     5 => B"00000001_000_0_1110",
     6 => B"000000000_000_0001",
     7 => B"00000000_000_1_1010",
     8 => B"00000000_000_0_0110",
     9 => B"00000000_110_0_1010",
     10 => B"000000000_000_1100",
     11 => B"00000000_101_1_1010",
     12 => B"00100000_000_0_1110",
     13 => B"000000000_101_0111",
     14 => B"10010_1110101_1101", 
     15 => B"00000000_010_1_1110",
     16 => B"00000010_001_1_1110",
     17 => B"00000010_000_0_1110",
     18 => B"000000000_001_0001",
     19 => B"00000000_001_1_1010",
     20 => B"00000000_010_0_1010",
     21 => B"00000000_001_0_0110",
     22 => B"00000000_110_0_1010",
     23 => B"000000000_001_1100",
     24 => B"00000000_101_1_1010",
     25 => B"00100000_000_0_1110",
     26 => B"000000000_101_0111",
     27 => B"10010_1110110_1101",
     28 => B"00000000_010_1_1110",
     29 => B"00000011_001_1_1110",
     30 => B"00000011_000_0_1110",
     31 => B"000000000_001_0001",
     32 => B"00000000_001_1_1010",
     33 => B"00000000_010_0_1010",
     34 => B"00000000_001_0_0110",
     35 => B"00000000_110_0_1010",
     36 => B"000000000_001_1100",
     37 => B"00000000_101_1_1010",
     38 => B"00100000_000_0_1110",
     39 => B"000000000_101_0111",
     40 => B"10010_1110110_1101",
     41 => B"00000000_010_1_1110",
     42 => B"00000101_001_1_1110",
     43 => B"00000101_000_0_1110",
     44 => B"000000000_001_0001",
     45 => B"00000000_001_1_1010",
     46 => B"00000000_010_0_1010",
     47 => B"00000000_001_0_0110",
     48 => B"00000000_110_0_1010",
     49 => B"000000000_001_1100",
     50 => B"00000000_101_1_1010",
     51 => B"00100000_000_0_1110",
     52 => B"000000000_101_0111",
     53 => B"10010_1110110_1101",
     54 => B"00000000_010_1_1110",
     55 => B"00000111_001_1_1110",
     56 => B"00000111_000_0_1110",
     57 => B"000000000_001_0001",
     58 => B"00000000_001_1_1010",
     59 => B"00000000_010_0_1010",
     60 => B"00000000_001_0_0110",
     61 => B"00000000_110_0_1010",
     62 => B"000000000_001_1100",
     63 => B"00000000_101_1_1010",
     64 => B"00100000_000_0_1110",
     65 => B"000000000_101_0111",
     66 => B"10010_1110110_1101",
     67 => B"00000000_010_1_1110",
     68 => B"00001011_001_1_1110",
     69 => B"00001011_000_0_1110",
     70 => B"000000000_001_0001",
     71 => B"00000000_001_1_1010",
     72 => B"00000000_010_0_1010",
     73 => B"00000000_001_0_0110",
     74 => B"00000000_110_0_1010",
     75 => B"000000000_001_1100",
     76 => B"00000000_101_1_1010",
     77 => B"00100000_000_0_1110",
     78 => B"000000000_101_0111",
     79 => B"10010_1110110_1101",
     80 => B"00000001_000_1_1110",
     81 => B"00000001_000_0_1110",
     82 => B"000000000_000_0001",
     83 => B"00000000_000_1_1010",
     84 => B"00000000_000_1_0110",
     85 => B"00000000_111_1_1010",
     86 => B"00100000_000_0_1110",
     87 => B"000000000_000_0111",
     88 => B"10010_1111001_1101",

       -- 0 => B"00000101_011_1_1110",
       -- 1 => B"00000000_100_1_1110",
       -- 2 => B"00000000_011_0_1010",
       -- 3 => B"000000000_100_0001",
       -- 4 => B"00000000_100_1_1010",
       -- 5 => B"00000001_000_0_1110",
       -- 6 => B"000000000_011_0001",
       -- 7 => B"00000000_011_1_1010",
       -- 8 => B"000011110_011_0100",
       -- 9 => B"00000_1111001_1101",
       -- 10 => B"00000000_100_0_1010",
       -- 11 => B"00000000_101_1_1010",

		others => (others => '0')
	);
	begin
		
	process(clk) begin
			
		if(rising_edge(clk)) then
			instout <= conteudo_rom(to_integer(address));
		end if;
	end process;
end architecture;	